.include gpdk90nm_ss.cir
.include param.cir
vdd 1 0 vdd_value
* --------------------------------------------------------------
* 2-Input NAND Gate
* Ports: inputA, inputB, Out, Vdd, Vss
* --------------------------------------------------------------
.subckt NAND_2 A B Out Vdd Vss

    * PMOS transistors
    XMP1 Out A Vdd Vdd pmos1v w=P_Width l=P_Length 
    XMP2 Out A Vdd Vdd pmos1v w=P_Width l=P_Length 

    * NMOS transistors
    XMN1 Out B N1 Vss nmos1v w=N_Width l=N_Length 
    XMN2 N1 B Vss Vss nmos1v w=N_Width l=N_Length 

.ends

* --------------------------------------------------------------
* 3-Input NAND Gate
* Ports: InputA, InputB, InputC, Output, Vdd, Vss
* --------------------------------------------------------------
.subckt NAND_3 A B Output Vdd Vss

    * PMOS transistors
    XMP1 Output A Vdd Vdd pmos1v w=P_Width l=P_Length 
    XMP2 Output A Vdd Vdd pmos1v w=P_Width l=P_Length
    XMP3 Output A Vdd Vdd pmos1v w=P_Width l=P_Length

    * NMOS transistors
    XMN1 Output B N1 Vss nmos1v w=N_Width l=N_Length 
    XMN2 N1 B N2 Vss nmos1v w=N_Width l=N_Length
    XMN3 N2 B Vss Vss nmos1v w=N_Width l=N_Length  

.ends
* --------------------------------------------------------------
* NAND Gates Implementation using PMOS and NMOS transistors
* --------------------------------------------------------------


* Instantiation of NAND gates
xNAND_2 1 0 out1 1 0 NAND_2
xNAND_3 1 0 out2 1 0 NAND_3

* --------------------------------------------------------------
* Simulation directives and plot commands
* --------------------------------------------------------------
.tran 0.0001n 2000n 500n

* Plots for NMOS current


.include DFFFF.cir
.option temp=00
.include waveW1.cir
.tran 0.001n 130n 100n
.plot v(Data) v(Clk) v(Out)
eW1.cir
.
*Waveform: 1100
vclk Clk 0 pulse    (vdd_value  0    5n     0.1n    0.1n    5000n     5001n)     
vd  Data 0 pulse    (0  vdd_value    5n     0.1n    0.1n    5000n     5001n)   
vres Reset 0 pulse  (0  vdd_value    5n     0.1n    0.1n    5000n     5001n)   
.tran 0.01 9000n 5100n
*Waveform 2: To Test the Datasampling when Data stays the same for a few Clock Edges
vclk Clk 0 pulse (0 vdd_value 5n 0.1n 0.1n 10n 20n)     
vres Reset 0 pulse (0 vdd_value 0 0.1n 0.1n 0n 0n)       
vd  Data 0 pulse (0 vdd_value 10n pRiseT pFallT 35n 80n) 
.tran 0.001n 200n 10n
